// SM_MCU.v

// Generated using ACDS version 14.0 200 at 2014.09.05.11:33:20

`timescale 1 ps / 1 ps
module SM_MCU (
		input  wire        clk_in_clk,          //       clk_in.clk
		input  wire        reset_in_reset_n,    //     reset_in.reset_n
		output wire [12:0] sdram_wire_addr,     //   sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,       //             .ba
		output wire        sdram_wire_cas_n,    //             .cas_n
		output wire        sdram_wire_cke,      //             .cke
		output wire        sdram_wire_cs_n,     //             .cs_n
		inout  wire [15:0] sdram_wire_dq,       //             .dq
		output wire [1:0]  sdram_wire_dqm,      //             .dqm
		output wire        sdram_wire_ras_n,    //             .ras_n
		output wire        sdram_wire_we_n,     //             .we_n
		output wire [1:0]  pio_led_export,      //      pio_led.export
		output wire [15:0] lcd_data_out_export, // lcd_data_out.export
		output wire        lcd_rs_export,       //       lcd_rs.export
		output wire        lcd_wr_export,       //       lcd_wr.export
		output wire        lcd_cs_export,       //       lcd_cs.export
		output wire        lcd_rd_export,       //       lcd_rd.export
		output wire        lcd_reset_export,    //    lcd_reset.export
		output wire        scl_export,          //          scl.export
		inout  wire        sda_export,          //          sda.export
		input  wire [1:0]  vs_int_in_export,    //    vs_int_in.export
		output wire        sm_2strobe_export,   //   sm_2strobe.export
		output wire        sm_1clr_export,      //      sm_1clr.export
		output wire        sm_1ena_export,      //      sm_1ena.export
		output wire [1:0]  sm_mux_export,       //       sm_mux.export
		input  wire [31:0] sm_data_in_export    //   sm_data_in.export
	);

	wire         cpu_instruction_master_waitrequest;                                // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                                    // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                                       // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                                   // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_readdatavalid;                              // mm_interconnect_0:CPU_instruction_master_readdatavalid -> CPU:i_readdatavalid
	wire         cpu_data_master_waitrequest;                                       // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                         // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [26:0] cpu_data_master_address;                                           // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire         cpu_data_master_write;                                             // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire         cpu_data_master_read;                                              // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                          // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_debugaccess;                                       // CPU:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire         cpu_data_master_readdatavalid;                                     // mm_interconnect_0:CPU_data_master_readdatavalid -> CPU:d_readdatavalid
	wire   [3:0] cpu_data_master_byteenable;                                        // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;               // CPU:jtag_debug_module_waitrequest -> mm_interconnect_0:CPU_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;                 // mm_interconnect_0:CPU_jtag_debug_module_writedata -> CPU:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                   // mm_interconnect_0:CPU_jtag_debug_module_address -> CPU:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                     // mm_interconnect_0:CPU_jtag_debug_module_write -> CPU:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                      // mm_interconnect_0:CPU_jtag_debug_module_read -> CPU:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                  // CPU:jtag_debug_module_readdata -> mm_interconnect_0:CPU_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;               // mm_interconnect_0:CPU_jtag_debug_module_debugaccess -> CPU:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;                // mm_interconnect_0:CPU_jtag_debug_module_byteenable -> CPU:jtag_debug_module_byteenable
	wire         mm_interconnect_0_sdram_s1_waitrequest;                            // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                              // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                                // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                             // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                                  // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                                   // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                               // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                          // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                             // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;         // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;            // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                            // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire   [1:0] mm_interconnect_0_pio_led_s1_address;                              // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_chipselect;                           // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire         mm_interconnect_0_pio_led_s1_write;                                // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                             // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;               // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                      // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire   [9:0] mm_interconnect_0_onchip_memory_s1_address;                        // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                     // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire         mm_interconnect_0_onchip_memory_s1_clken;                          // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_onchip_memory_s1_write;                          // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                       // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                     // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire  [31:0] mm_interconnect_0_lcd_data_out_s1_writedata;                       // mm_interconnect_0:LCD_DATA_OUT_s1_writedata -> LCD_DATA_OUT:writedata
	wire   [1:0] mm_interconnect_0_lcd_data_out_s1_address;                         // mm_interconnect_0:LCD_DATA_OUT_s1_address -> LCD_DATA_OUT:address
	wire         mm_interconnect_0_lcd_data_out_s1_chipselect;                      // mm_interconnect_0:LCD_DATA_OUT_s1_chipselect -> LCD_DATA_OUT:chipselect
	wire         mm_interconnect_0_lcd_data_out_s1_write;                           // mm_interconnect_0:LCD_DATA_OUT_s1_write -> LCD_DATA_OUT:write_n
	wire  [31:0] mm_interconnect_0_lcd_data_out_s1_readdata;                        // LCD_DATA_OUT:readdata -> mm_interconnect_0:LCD_DATA_OUT_s1_readdata
	wire  [31:0] mm_interconnect_0_lcd_rs_s1_writedata;                             // mm_interconnect_0:LCD_RS_s1_writedata -> LCD_RS:writedata
	wire   [1:0] mm_interconnect_0_lcd_rs_s1_address;                               // mm_interconnect_0:LCD_RS_s1_address -> LCD_RS:address
	wire         mm_interconnect_0_lcd_rs_s1_chipselect;                            // mm_interconnect_0:LCD_RS_s1_chipselect -> LCD_RS:chipselect
	wire         mm_interconnect_0_lcd_rs_s1_write;                                 // mm_interconnect_0:LCD_RS_s1_write -> LCD_RS:write_n
	wire  [31:0] mm_interconnect_0_lcd_rs_s1_readdata;                              // LCD_RS:readdata -> mm_interconnect_0:LCD_RS_s1_readdata
	wire  [31:0] mm_interconnect_0_lcd_wr_s1_writedata;                             // mm_interconnect_0:LCD_WR_s1_writedata -> LCD_WR:writedata
	wire   [1:0] mm_interconnect_0_lcd_wr_s1_address;                               // mm_interconnect_0:LCD_WR_s1_address -> LCD_WR:address
	wire         mm_interconnect_0_lcd_wr_s1_chipselect;                            // mm_interconnect_0:LCD_WR_s1_chipselect -> LCD_WR:chipselect
	wire         mm_interconnect_0_lcd_wr_s1_write;                                 // mm_interconnect_0:LCD_WR_s1_write -> LCD_WR:write_n
	wire  [31:0] mm_interconnect_0_lcd_wr_s1_readdata;                              // LCD_WR:readdata -> mm_interconnect_0:LCD_WR_s1_readdata
	wire  [31:0] mm_interconnect_0_lcd_cs_s1_writedata;                             // mm_interconnect_0:LCD_CS_s1_writedata -> LCD_CS:writedata
	wire   [1:0] mm_interconnect_0_lcd_cs_s1_address;                               // mm_interconnect_0:LCD_CS_s1_address -> LCD_CS:address
	wire         mm_interconnect_0_lcd_cs_s1_chipselect;                            // mm_interconnect_0:LCD_CS_s1_chipselect -> LCD_CS:chipselect
	wire         mm_interconnect_0_lcd_cs_s1_write;                                 // mm_interconnect_0:LCD_CS_s1_write -> LCD_CS:write_n
	wire  [31:0] mm_interconnect_0_lcd_cs_s1_readdata;                              // LCD_CS:readdata -> mm_interconnect_0:LCD_CS_s1_readdata
	wire  [31:0] mm_interconnect_0_lcd_reset_s1_writedata;                          // mm_interconnect_0:LCD_RESET_s1_writedata -> LCD_RESET:writedata
	wire   [1:0] mm_interconnect_0_lcd_reset_s1_address;                            // mm_interconnect_0:LCD_RESET_s1_address -> LCD_RESET:address
	wire         mm_interconnect_0_lcd_reset_s1_chipselect;                         // mm_interconnect_0:LCD_RESET_s1_chipselect -> LCD_RESET:chipselect
	wire         mm_interconnect_0_lcd_reset_s1_write;                              // mm_interconnect_0:LCD_RESET_s1_write -> LCD_RESET:write_n
	wire  [31:0] mm_interconnect_0_lcd_reset_s1_readdata;                           // LCD_RESET:readdata -> mm_interconnect_0:LCD_RESET_s1_readdata
	wire  [31:0] mm_interconnect_0_sda_s1_writedata;                                // mm_interconnect_0:SDA_s1_writedata -> SDA:writedata
	wire   [1:0] mm_interconnect_0_sda_s1_address;                                  // mm_interconnect_0:SDA_s1_address -> SDA:address
	wire         mm_interconnect_0_sda_s1_chipselect;                               // mm_interconnect_0:SDA_s1_chipselect -> SDA:chipselect
	wire         mm_interconnect_0_sda_s1_write;                                    // mm_interconnect_0:SDA_s1_write -> SDA:write_n
	wire  [31:0] mm_interconnect_0_sda_s1_readdata;                                 // SDA:readdata -> mm_interconnect_0:SDA_s1_readdata
	wire  [31:0] mm_interconnect_0_sm_1clr_s1_writedata;                            // mm_interconnect_0:SM_1clr_s1_writedata -> SM_1clr:writedata
	wire   [1:0] mm_interconnect_0_sm_1clr_s1_address;                              // mm_interconnect_0:SM_1clr_s1_address -> SM_1clr:address
	wire         mm_interconnect_0_sm_1clr_s1_chipselect;                           // mm_interconnect_0:SM_1clr_s1_chipselect -> SM_1clr:chipselect
	wire         mm_interconnect_0_sm_1clr_s1_write;                                // mm_interconnect_0:SM_1clr_s1_write -> SM_1clr:write_n
	wire  [31:0] mm_interconnect_0_sm_1clr_s1_readdata;                             // SM_1clr:readdata -> mm_interconnect_0:SM_1clr_s1_readdata
	wire  [31:0] mm_interconnect_0_sm_1ena_s1_writedata;                            // mm_interconnect_0:SM_1ena_s1_writedata -> SM_1ena:writedata
	wire   [1:0] mm_interconnect_0_sm_1ena_s1_address;                              // mm_interconnect_0:SM_1ena_s1_address -> SM_1ena:address
	wire         mm_interconnect_0_sm_1ena_s1_chipselect;                           // mm_interconnect_0:SM_1ena_s1_chipselect -> SM_1ena:chipselect
	wire         mm_interconnect_0_sm_1ena_s1_write;                                // mm_interconnect_0:SM_1ena_s1_write -> SM_1ena:write_n
	wire  [31:0] mm_interconnect_0_sm_1ena_s1_readdata;                             // SM_1ena:readdata -> mm_interconnect_0:SM_1ena_s1_readdata
	wire  [31:0] mm_interconnect_0_sm_mux_s1_writedata;                             // mm_interconnect_0:SM_mux_s1_writedata -> SM_mux:writedata
	wire   [1:0] mm_interconnect_0_sm_mux_s1_address;                               // mm_interconnect_0:SM_mux_s1_address -> SM_mux:address
	wire         mm_interconnect_0_sm_mux_s1_chipselect;                            // mm_interconnect_0:SM_mux_s1_chipselect -> SM_mux:chipselect
	wire         mm_interconnect_0_sm_mux_s1_write;                                 // mm_interconnect_0:SM_mux_s1_write -> SM_mux:write_n
	wire  [31:0] mm_interconnect_0_sm_mux_s1_readdata;                              // SM_mux:readdata -> mm_interconnect_0:SM_mux_s1_readdata
	wire   [1:0] mm_interconnect_0_sm_data_in_s1_address;                           // mm_interconnect_0:SM_data_in_s1_address -> SM_data_in:address
	wire  [31:0] mm_interconnect_0_sm_data_in_s1_readdata;                          // SM_data_in:readdata -> mm_interconnect_0:SM_data_in_s1_readdata
	wire  [31:0] mm_interconnect_0_lcd_rd_s1_writedata;                             // mm_interconnect_0:LCD_RD_s1_writedata -> LCD_RD:writedata
	wire   [1:0] mm_interconnect_0_lcd_rd_s1_address;                               // mm_interconnect_0:LCD_RD_s1_address -> LCD_RD:address
	wire         mm_interconnect_0_lcd_rd_s1_chipselect;                            // mm_interconnect_0:LCD_RD_s1_chipselect -> LCD_RD:chipselect
	wire         mm_interconnect_0_lcd_rd_s1_write;                                 // mm_interconnect_0:LCD_RD_s1_write -> LCD_RD:write_n
	wire  [31:0] mm_interconnect_0_lcd_rd_s1_readdata;                              // LCD_RD:readdata -> mm_interconnect_0:LCD_RD_s1_readdata
	wire  [31:0] mm_interconnect_0_vs_int_in_s1_writedata;                          // mm_interconnect_0:VS_int_in_s1_writedata -> VS_int_in:writedata
	wire   [1:0] mm_interconnect_0_vs_int_in_s1_address;                            // mm_interconnect_0:VS_int_in_s1_address -> VS_int_in:address
	wire         mm_interconnect_0_vs_int_in_s1_chipselect;                         // mm_interconnect_0:VS_int_in_s1_chipselect -> VS_int_in:chipselect
	wire         mm_interconnect_0_vs_int_in_s1_write;                              // mm_interconnect_0:VS_int_in_s1_write -> VS_int_in:write_n
	wire  [31:0] mm_interconnect_0_vs_int_in_s1_readdata;                           // VS_int_in:readdata -> mm_interconnect_0:VS_int_in_s1_readdata
	wire  [31:0] mm_interconnect_0_performance_counter_control_slave_writedata;     // mm_interconnect_0:performance_counter_control_slave_writedata -> performance_counter:writedata
	wire   [3:0] mm_interconnect_0_performance_counter_control_slave_address;       // mm_interconnect_0:performance_counter_control_slave_address -> performance_counter:address
	wire         mm_interconnect_0_performance_counter_control_slave_write;         // mm_interconnect_0:performance_counter_control_slave_write -> performance_counter:write
	wire  [31:0] mm_interconnect_0_performance_counter_control_slave_readdata;      // performance_counter:readdata -> mm_interconnect_0:performance_counter_control_slave_readdata
	wire         mm_interconnect_0_performance_counter_control_slave_begintransfer; // mm_interconnect_0:performance_counter_control_slave_begintransfer -> performance_counter:begintransfer
	wire  [31:0] mm_interconnect_0_sm_2strobe_s1_writedata;                         // mm_interconnect_0:SM_2strobe_s1_writedata -> SM_2strobe:writedata
	wire   [1:0] mm_interconnect_0_sm_2strobe_s1_address;                           // mm_interconnect_0:SM_2strobe_s1_address -> SM_2strobe:address
	wire         mm_interconnect_0_sm_2strobe_s1_chipselect;                        // mm_interconnect_0:SM_2strobe_s1_chipselect -> SM_2strobe:chipselect
	wire         mm_interconnect_0_sm_2strobe_s1_write;                             // mm_interconnect_0:SM_2strobe_s1_write -> SM_2strobe:write_n
	wire  [31:0] mm_interconnect_0_sm_2strobe_s1_readdata;                          // SM_2strobe:readdata -> mm_interconnect_0:SM_2strobe_s1_readdata
	wire  [31:0] mm_interconnect_0_scl_s1_writedata;                                // mm_interconnect_0:SCL_s1_writedata -> SCL:writedata
	wire   [1:0] mm_interconnect_0_scl_s1_address;                                  // mm_interconnect_0:SCL_s1_address -> SCL:address
	wire         mm_interconnect_0_scl_s1_chipselect;                               // mm_interconnect_0:SCL_s1_chipselect -> SCL:chipselect
	wire         mm_interconnect_0_scl_s1_write;                                    // mm_interconnect_0:SCL_s1_write -> SCL:write_n
	wire  [31:0] mm_interconnect_0_scl_s1_readdata;                                 // SCL:readdata -> mm_interconnect_0:SCL_s1_readdata
	wire         irq_mapper_receiver0_irq;                                          // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                          // VS_int_in:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_d_irq_irq;                                                     // irq_mapper:sender_irq -> CPU:d_irq
	wire         rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [CPU:reset_n, LCD_CS:reset_n, LCD_DATA_OUT:reset_n, LCD_RD:reset_n, LCD_RESET:reset_n, LCD_RS:reset_n, LCD_WR:reset_n, SCL:reset_n, SDA:reset_n, SM_1clr:reset_n, SM_1ena:reset_n, SM_2strobe:reset_n, SM_data_in:reset_n, SM_mux:reset_n, VS_int_in:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:CPU_reset_n_reset_bridge_in_reset_reset, onchip_memory:reset, performance_counter:reset_n, pio_led:reset_n, rst_translator:in_reset, sdram:reset_n, sysid_qsys:reset_n]
	wire         rst_controller_reset_out_reset_req;                                // rst_controller:reset_req -> [CPU:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                                 // CPU:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	SM_MCU_sdram sdram (
		.clk            (clk_in_clk),                               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	SM_MCU_pio_led pio_led (
		.clk        (clk_in_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_export)                           // external_connection.export
	);

	SM_MCU_jtag_uart jtag_uart (
		.clk            (clk_in_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	SM_MCU_onchip_memory onchip_memory (
		.clk        (clk_in_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	SM_MCU_LCD_DATA_OUT lcd_data_out (
		.clk        (clk_in_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_lcd_data_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_data_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_data_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_data_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_data_out_s1_readdata),   //                    .readdata
		.out_port   (lcd_data_out_export)                           // external_connection.export
	);

	SM_MCU_LCD_RS lcd_rs (
		.clk        (clk_in_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_lcd_rs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_rs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_rs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_rs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_rs_s1_readdata),   //                    .readdata
		.out_port   (lcd_rs_export)                           // external_connection.export
	);

	SM_MCU_LCD_RS lcd_wr (
		.clk        (clk_in_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_lcd_wr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_wr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_wr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_wr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_wr_s1_readdata),   //                    .readdata
		.out_port   (lcd_wr_export)                           // external_connection.export
	);

	SM_MCU_LCD_RS lcd_rd (
		.clk        (clk_in_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_lcd_rd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_rd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_rd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_rd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_rd_s1_readdata),   //                    .readdata
		.out_port   (lcd_rd_export)                           // external_connection.export
	);

	SM_MCU_LCD_RS lcd_cs (
		.clk        (clk_in_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_lcd_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_cs_s1_readdata),   //                    .readdata
		.out_port   (lcd_cs_export)                           // external_connection.export
	);

	SM_MCU_LCD_RS lcd_reset (
		.clk        (clk_in_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_lcd_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_reset_s1_readdata),   //                    .readdata
		.out_port   (lcd_reset_export)                           // external_connection.export
	);

	SM_MCU_SCL scl (
		.clk        (clk_in_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_scl_s1_readdata),   //                    .readdata
		.out_port   (scl_export)                           // external_connection.export
	);

	SM_MCU_SDA sda (
		.clk        (clk_in_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sda_s1_readdata),   //                    .readdata
		.bidir_port (sda_export)                           // external_connection.export
	);

	SM_MCU_performance_counter performance_counter (
		.clk           (clk_in_clk),                                                        //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                   //         reset.reset_n
		.address       (mm_interconnect_0_performance_counter_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_0_performance_counter_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_0_performance_counter_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_0_performance_counter_control_slave_write),         //              .write
		.writedata     (mm_interconnect_0_performance_counter_control_slave_writedata)      //              .writedata
	);

	SM_MCU_CPU cpu (
		.clk                                   (clk_in_clk),                                          //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	SM_MCU_sysid_qsys sysid_qsys (
		.clock    (clk_in_clk),                                          //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	SM_MCU_VS_int_in vs_int_in (
		.clk        (clk_in_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_vs_int_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_vs_int_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_vs_int_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_vs_int_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_vs_int_in_s1_readdata),   //                    .readdata
		.in_port    (vs_int_in_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                   //                 irq.irq
	);

	SM_MCU_LCD_RS sm_2strobe (
		.clk        (clk_in_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_sm_2strobe_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sm_2strobe_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sm_2strobe_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sm_2strobe_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sm_2strobe_s1_readdata),   //                    .readdata
		.out_port   (sm_2strobe_export)                           // external_connection.export
	);

	SM_MCU_SCL sm_1clr (
		.clk        (clk_in_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_sm_1clr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sm_1clr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sm_1clr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sm_1clr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sm_1clr_s1_readdata),   //                    .readdata
		.out_port   (sm_1clr_export)                           // external_connection.export
	);

	SM_MCU_LCD_RS sm_1ena (
		.clk        (clk_in_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_sm_1ena_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sm_1ena_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sm_1ena_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sm_1ena_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sm_1ena_s1_readdata),   //                    .readdata
		.out_port   (sm_1ena_export)                           // external_connection.export
	);

	SM_MCU_SM_mux sm_mux (
		.clk        (clk_in_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_sm_mux_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sm_mux_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sm_mux_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sm_mux_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sm_mux_s1_readdata),   //                    .readdata
		.out_port   (sm_mux_export)                           // external_connection.export
	);

	SM_MCU_SM_data_in sm_data_in (
		.clk      (clk_in_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_sm_data_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sm_data_in_s1_readdata), //                    .readdata
		.in_port  (sm_data_in_export)                         // external_connection.export
	);

	SM_MCU_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                     (clk_in_clk),                                                        //                           clk_clk.clk
		.CPU_reset_n_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                                    // CPU_reset_n_reset_bridge_in_reset.reset
		.CPU_data_master_address                         (cpu_data_master_address),                                           //                   CPU_data_master.address
		.CPU_data_master_waitrequest                     (cpu_data_master_waitrequest),                                       //                                  .waitrequest
		.CPU_data_master_byteenable                      (cpu_data_master_byteenable),                                        //                                  .byteenable
		.CPU_data_master_read                            (cpu_data_master_read),                                              //                                  .read
		.CPU_data_master_readdata                        (cpu_data_master_readdata),                                          //                                  .readdata
		.CPU_data_master_readdatavalid                   (cpu_data_master_readdatavalid),                                     //                                  .readdatavalid
		.CPU_data_master_write                           (cpu_data_master_write),                                             //                                  .write
		.CPU_data_master_writedata                       (cpu_data_master_writedata),                                         //                                  .writedata
		.CPU_data_master_debugaccess                     (cpu_data_master_debugaccess),                                       //                                  .debugaccess
		.CPU_instruction_master_address                  (cpu_instruction_master_address),                                    //            CPU_instruction_master.address
		.CPU_instruction_master_waitrequest              (cpu_instruction_master_waitrequest),                                //                                  .waitrequest
		.CPU_instruction_master_read                     (cpu_instruction_master_read),                                       //                                  .read
		.CPU_instruction_master_readdata                 (cpu_instruction_master_readdata),                                   //                                  .readdata
		.CPU_instruction_master_readdatavalid            (cpu_instruction_master_readdatavalid),                              //                                  .readdatavalid
		.CPU_jtag_debug_module_address                   (mm_interconnect_0_cpu_jtag_debug_module_address),                   //             CPU_jtag_debug_module.address
		.CPU_jtag_debug_module_write                     (mm_interconnect_0_cpu_jtag_debug_module_write),                     //                                  .write
		.CPU_jtag_debug_module_read                      (mm_interconnect_0_cpu_jtag_debug_module_read),                      //                                  .read
		.CPU_jtag_debug_module_readdata                  (mm_interconnect_0_cpu_jtag_debug_module_readdata),                  //                                  .readdata
		.CPU_jtag_debug_module_writedata                 (mm_interconnect_0_cpu_jtag_debug_module_writedata),                 //                                  .writedata
		.CPU_jtag_debug_module_byteenable                (mm_interconnect_0_cpu_jtag_debug_module_byteenable),                //                                  .byteenable
		.CPU_jtag_debug_module_waitrequest               (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),               //                                  .waitrequest
		.CPU_jtag_debug_module_debugaccess               (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),               //                                  .debugaccess
		.jtag_uart_avalon_jtag_slave_address             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),             //       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),               //                                  .write
		.jtag_uart_avalon_jtag_slave_read                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                //                                  .read
		.jtag_uart_avalon_jtag_slave_readdata            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),            //                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),           //                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),         //                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),          //                                  .chipselect
		.LCD_CS_s1_address                               (mm_interconnect_0_lcd_cs_s1_address),                               //                         LCD_CS_s1.address
		.LCD_CS_s1_write                                 (mm_interconnect_0_lcd_cs_s1_write),                                 //                                  .write
		.LCD_CS_s1_readdata                              (mm_interconnect_0_lcd_cs_s1_readdata),                              //                                  .readdata
		.LCD_CS_s1_writedata                             (mm_interconnect_0_lcd_cs_s1_writedata),                             //                                  .writedata
		.LCD_CS_s1_chipselect                            (mm_interconnect_0_lcd_cs_s1_chipselect),                            //                                  .chipselect
		.LCD_DATA_OUT_s1_address                         (mm_interconnect_0_lcd_data_out_s1_address),                         //                   LCD_DATA_OUT_s1.address
		.LCD_DATA_OUT_s1_write                           (mm_interconnect_0_lcd_data_out_s1_write),                           //                                  .write
		.LCD_DATA_OUT_s1_readdata                        (mm_interconnect_0_lcd_data_out_s1_readdata),                        //                                  .readdata
		.LCD_DATA_OUT_s1_writedata                       (mm_interconnect_0_lcd_data_out_s1_writedata),                       //                                  .writedata
		.LCD_DATA_OUT_s1_chipselect                      (mm_interconnect_0_lcd_data_out_s1_chipselect),                      //                                  .chipselect
		.LCD_RD_s1_address                               (mm_interconnect_0_lcd_rd_s1_address),                               //                         LCD_RD_s1.address
		.LCD_RD_s1_write                                 (mm_interconnect_0_lcd_rd_s1_write),                                 //                                  .write
		.LCD_RD_s1_readdata                              (mm_interconnect_0_lcd_rd_s1_readdata),                              //                                  .readdata
		.LCD_RD_s1_writedata                             (mm_interconnect_0_lcd_rd_s1_writedata),                             //                                  .writedata
		.LCD_RD_s1_chipselect                            (mm_interconnect_0_lcd_rd_s1_chipselect),                            //                                  .chipselect
		.LCD_RESET_s1_address                            (mm_interconnect_0_lcd_reset_s1_address),                            //                      LCD_RESET_s1.address
		.LCD_RESET_s1_write                              (mm_interconnect_0_lcd_reset_s1_write),                              //                                  .write
		.LCD_RESET_s1_readdata                           (mm_interconnect_0_lcd_reset_s1_readdata),                           //                                  .readdata
		.LCD_RESET_s1_writedata                          (mm_interconnect_0_lcd_reset_s1_writedata),                          //                                  .writedata
		.LCD_RESET_s1_chipselect                         (mm_interconnect_0_lcd_reset_s1_chipselect),                         //                                  .chipselect
		.LCD_RS_s1_address                               (mm_interconnect_0_lcd_rs_s1_address),                               //                         LCD_RS_s1.address
		.LCD_RS_s1_write                                 (mm_interconnect_0_lcd_rs_s1_write),                                 //                                  .write
		.LCD_RS_s1_readdata                              (mm_interconnect_0_lcd_rs_s1_readdata),                              //                                  .readdata
		.LCD_RS_s1_writedata                             (mm_interconnect_0_lcd_rs_s1_writedata),                             //                                  .writedata
		.LCD_RS_s1_chipselect                            (mm_interconnect_0_lcd_rs_s1_chipselect),                            //                                  .chipselect
		.LCD_WR_s1_address                               (mm_interconnect_0_lcd_wr_s1_address),                               //                         LCD_WR_s1.address
		.LCD_WR_s1_write                                 (mm_interconnect_0_lcd_wr_s1_write),                                 //                                  .write
		.LCD_WR_s1_readdata                              (mm_interconnect_0_lcd_wr_s1_readdata),                              //                                  .readdata
		.LCD_WR_s1_writedata                             (mm_interconnect_0_lcd_wr_s1_writedata),                             //                                  .writedata
		.LCD_WR_s1_chipselect                            (mm_interconnect_0_lcd_wr_s1_chipselect),                            //                                  .chipselect
		.onchip_memory_s1_address                        (mm_interconnect_0_onchip_memory_s1_address),                        //                  onchip_memory_s1.address
		.onchip_memory_s1_write                          (mm_interconnect_0_onchip_memory_s1_write),                          //                                  .write
		.onchip_memory_s1_readdata                       (mm_interconnect_0_onchip_memory_s1_readdata),                       //                                  .readdata
		.onchip_memory_s1_writedata                      (mm_interconnect_0_onchip_memory_s1_writedata),                      //                                  .writedata
		.onchip_memory_s1_byteenable                     (mm_interconnect_0_onchip_memory_s1_byteenable),                     //                                  .byteenable
		.onchip_memory_s1_chipselect                     (mm_interconnect_0_onchip_memory_s1_chipselect),                     //                                  .chipselect
		.onchip_memory_s1_clken                          (mm_interconnect_0_onchip_memory_s1_clken),                          //                                  .clken
		.performance_counter_control_slave_address       (mm_interconnect_0_performance_counter_control_slave_address),       // performance_counter_control_slave.address
		.performance_counter_control_slave_write         (mm_interconnect_0_performance_counter_control_slave_write),         //                                  .write
		.performance_counter_control_slave_readdata      (mm_interconnect_0_performance_counter_control_slave_readdata),      //                                  .readdata
		.performance_counter_control_slave_writedata     (mm_interconnect_0_performance_counter_control_slave_writedata),     //                                  .writedata
		.performance_counter_control_slave_begintransfer (mm_interconnect_0_performance_counter_control_slave_begintransfer), //                                  .begintransfer
		.pio_led_s1_address                              (mm_interconnect_0_pio_led_s1_address),                              //                        pio_led_s1.address
		.pio_led_s1_write                                (mm_interconnect_0_pio_led_s1_write),                                //                                  .write
		.pio_led_s1_readdata                             (mm_interconnect_0_pio_led_s1_readdata),                             //                                  .readdata
		.pio_led_s1_writedata                            (mm_interconnect_0_pio_led_s1_writedata),                            //                                  .writedata
		.pio_led_s1_chipselect                           (mm_interconnect_0_pio_led_s1_chipselect),                           //                                  .chipselect
		.SCL_s1_address                                  (mm_interconnect_0_scl_s1_address),                                  //                            SCL_s1.address
		.SCL_s1_write                                    (mm_interconnect_0_scl_s1_write),                                    //                                  .write
		.SCL_s1_readdata                                 (mm_interconnect_0_scl_s1_readdata),                                 //                                  .readdata
		.SCL_s1_writedata                                (mm_interconnect_0_scl_s1_writedata),                                //                                  .writedata
		.SCL_s1_chipselect                               (mm_interconnect_0_scl_s1_chipselect),                               //                                  .chipselect
		.SDA_s1_address                                  (mm_interconnect_0_sda_s1_address),                                  //                            SDA_s1.address
		.SDA_s1_write                                    (mm_interconnect_0_sda_s1_write),                                    //                                  .write
		.SDA_s1_readdata                                 (mm_interconnect_0_sda_s1_readdata),                                 //                                  .readdata
		.SDA_s1_writedata                                (mm_interconnect_0_sda_s1_writedata),                                //                                  .writedata
		.SDA_s1_chipselect                               (mm_interconnect_0_sda_s1_chipselect),                               //                                  .chipselect
		.sdram_s1_address                                (mm_interconnect_0_sdram_s1_address),                                //                          sdram_s1.address
		.sdram_s1_write                                  (mm_interconnect_0_sdram_s1_write),                                  //                                  .write
		.sdram_s1_read                                   (mm_interconnect_0_sdram_s1_read),                                   //                                  .read
		.sdram_s1_readdata                               (mm_interconnect_0_sdram_s1_readdata),                               //                                  .readdata
		.sdram_s1_writedata                              (mm_interconnect_0_sdram_s1_writedata),                              //                                  .writedata
		.sdram_s1_byteenable                             (mm_interconnect_0_sdram_s1_byteenable),                             //                                  .byteenable
		.sdram_s1_readdatavalid                          (mm_interconnect_0_sdram_s1_readdatavalid),                          //                                  .readdatavalid
		.sdram_s1_waitrequest                            (mm_interconnect_0_sdram_s1_waitrequest),                            //                                  .waitrequest
		.sdram_s1_chipselect                             (mm_interconnect_0_sdram_s1_chipselect),                             //                                  .chipselect
		.SM_1clr_s1_address                              (mm_interconnect_0_sm_1clr_s1_address),                              //                        SM_1clr_s1.address
		.SM_1clr_s1_write                                (mm_interconnect_0_sm_1clr_s1_write),                                //                                  .write
		.SM_1clr_s1_readdata                             (mm_interconnect_0_sm_1clr_s1_readdata),                             //                                  .readdata
		.SM_1clr_s1_writedata                            (mm_interconnect_0_sm_1clr_s1_writedata),                            //                                  .writedata
		.SM_1clr_s1_chipselect                           (mm_interconnect_0_sm_1clr_s1_chipselect),                           //                                  .chipselect
		.SM_1ena_s1_address                              (mm_interconnect_0_sm_1ena_s1_address),                              //                        SM_1ena_s1.address
		.SM_1ena_s1_write                                (mm_interconnect_0_sm_1ena_s1_write),                                //                                  .write
		.SM_1ena_s1_readdata                             (mm_interconnect_0_sm_1ena_s1_readdata),                             //                                  .readdata
		.SM_1ena_s1_writedata                            (mm_interconnect_0_sm_1ena_s1_writedata),                            //                                  .writedata
		.SM_1ena_s1_chipselect                           (mm_interconnect_0_sm_1ena_s1_chipselect),                           //                                  .chipselect
		.SM_2strobe_s1_address                           (mm_interconnect_0_sm_2strobe_s1_address),                           //                     SM_2strobe_s1.address
		.SM_2strobe_s1_write                             (mm_interconnect_0_sm_2strobe_s1_write),                             //                                  .write
		.SM_2strobe_s1_readdata                          (mm_interconnect_0_sm_2strobe_s1_readdata),                          //                                  .readdata
		.SM_2strobe_s1_writedata                         (mm_interconnect_0_sm_2strobe_s1_writedata),                         //                                  .writedata
		.SM_2strobe_s1_chipselect                        (mm_interconnect_0_sm_2strobe_s1_chipselect),                        //                                  .chipselect
		.SM_data_in_s1_address                           (mm_interconnect_0_sm_data_in_s1_address),                           //                     SM_data_in_s1.address
		.SM_data_in_s1_readdata                          (mm_interconnect_0_sm_data_in_s1_readdata),                          //                                  .readdata
		.SM_mux_s1_address                               (mm_interconnect_0_sm_mux_s1_address),                               //                         SM_mux_s1.address
		.SM_mux_s1_write                                 (mm_interconnect_0_sm_mux_s1_write),                                 //                                  .write
		.SM_mux_s1_readdata                              (mm_interconnect_0_sm_mux_s1_readdata),                              //                                  .readdata
		.SM_mux_s1_writedata                             (mm_interconnect_0_sm_mux_s1_writedata),                             //                                  .writedata
		.SM_mux_s1_chipselect                            (mm_interconnect_0_sm_mux_s1_chipselect),                            //                                  .chipselect
		.sysid_qsys_control_slave_address                (mm_interconnect_0_sysid_qsys_control_slave_address),                //          sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata               (mm_interconnect_0_sysid_qsys_control_slave_readdata),               //                                  .readdata
		.VS_int_in_s1_address                            (mm_interconnect_0_vs_int_in_s1_address),                            //                      VS_int_in_s1.address
		.VS_int_in_s1_write                              (mm_interconnect_0_vs_int_in_s1_write),                              //                                  .write
		.VS_int_in_s1_readdata                           (mm_interconnect_0_vs_int_in_s1_readdata),                           //                                  .readdata
		.VS_int_in_s1_writedata                          (mm_interconnect_0_vs_int_in_s1_writedata),                          //                                  .writedata
		.VS_int_in_s1_chipselect                         (mm_interconnect_0_vs_int_in_s1_chipselect)                          //                                  .chipselect
	);

	SM_MCU_irq_mapper irq_mapper (
		.clk           (clk_in_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_in_reset_n),                  // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_in_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
